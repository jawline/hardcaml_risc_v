module op (
    funct7,
    rhs,
    lhs,
    funct3,
    new_rd,
    error
);

    input [6:0] funct7;
    input [31:0] rhs;
    input [31:0] lhs;
    input [2:0] funct3;
    output [31:0] new_rd;
    output error;

    /* signal declarations */
    wire _19 = 1'b0;
    wire _18 = 1'b0;
    wire [6:0] _16 = 7'b0000001;
    wire _17;
    wire _15 = 1'b0;
    wire _14 = 1'b0;
    wire _13 = 1'b0;
    wire _12 = 1'b0;
    wire _11 = 1'b0;
    reg _20;
    wire [31:0] _481;
    wire [31:0] _480;
    wire [31:0] _477 = 32'b11111111111111111111111111111111;
    wire _474;
    wire [2:0] _470;
    wire [6:0] _471;
    wire [14:0] _472;
    wire _465;
    wire [1:0] _466;
    wire [3:0] _467;
    wire [7:0] _468;
    wire [15:0] _469;
    wire [30:0] _473;
    wire [31:0] _475;
    wire [1:0] _463;
    wire [5:0] _460;
    wire [13:0] _461;
    wire _455;
    wire [1:0] _456;
    wire [3:0] _457;
    wire [7:0] _458;
    wire [15:0] _459;
    wire [29:0] _462;
    wire [31:0] _464;
    wire [2:0] _453;
    wire [4:0] _450;
    wire [12:0] _451;
    wire _445;
    wire [1:0] _446;
    wire [3:0] _447;
    wire [7:0] _448;
    wire [15:0] _449;
    wire [28:0] _452;
    wire [31:0] _454;
    wire [3:0] _443;
    wire [11:0] _441;
    wire _436;
    wire [1:0] _437;
    wire [3:0] _438;
    wire [7:0] _439;
    wire [15:0] _440;
    wire [27:0] _442;
    wire [31:0] _444;
    wire [4:0] _434;
    wire [2:0] _431;
    wire [10:0] _432;
    wire _426;
    wire [1:0] _427;
    wire [3:0] _428;
    wire [7:0] _429;
    wire [15:0] _430;
    wire [26:0] _433;
    wire [31:0] _435;
    wire [5:0] _424;
    wire [9:0] _422;
    wire _417;
    wire [1:0] _418;
    wire [3:0] _419;
    wire [7:0] _420;
    wire [15:0] _421;
    wire [25:0] _423;
    wire [31:0] _425;
    wire [6:0] _415;
    wire [8:0] _413;
    wire _408;
    wire [1:0] _409;
    wire [3:0] _410;
    wire [7:0] _411;
    wire [15:0] _412;
    wire [24:0] _414;
    wire [31:0] _416;
    wire [7:0] _406;
    wire _400;
    wire [1:0] _401;
    wire [3:0] _402;
    wire [7:0] _403;
    wire [15:0] _404;
    wire [23:0] _405;
    wire [31:0] _407;
    wire [8:0] _398;
    wire [2:0] _395;
    wire [6:0] _396;
    wire _390;
    wire [1:0] _391;
    wire [3:0] _392;
    wire [7:0] _393;
    wire [15:0] _394;
    wire [22:0] _397;
    wire [31:0] _399;
    wire [9:0] _388;
    wire [5:0] _386;
    wire _381;
    wire [1:0] _382;
    wire [3:0] _383;
    wire [7:0] _384;
    wire [15:0] _385;
    wire [21:0] _387;
    wire [31:0] _389;
    wire [10:0] _379;
    wire [4:0] _377;
    wire _372;
    wire [1:0] _373;
    wire [3:0] _374;
    wire [7:0] _375;
    wire [15:0] _376;
    wire [20:0] _378;
    wire [31:0] _380;
    wire [11:0] _370;
    wire _364;
    wire [1:0] _365;
    wire [3:0] _366;
    wire [7:0] _367;
    wire [15:0] _368;
    wire [19:0] _369;
    wire [31:0] _371;
    wire [12:0] _362;
    wire [2:0] _360;
    wire _355;
    wire [1:0] _356;
    wire [3:0] _357;
    wire [7:0] _358;
    wire [15:0] _359;
    wire [18:0] _361;
    wire [31:0] _363;
    wire [13:0] _353;
    wire _347;
    wire [1:0] _348;
    wire [3:0] _349;
    wire [7:0] _350;
    wire [15:0] _351;
    wire [17:0] _352;
    wire [31:0] _354;
    wire [14:0] _345;
    wire _339;
    wire [1:0] _340;
    wire [3:0] _341;
    wire [7:0] _342;
    wire [15:0] _343;
    wire [16:0] _344;
    wire [31:0] _346;
    wire [15:0] _337;
    wire _332;
    wire [1:0] _333;
    wire [3:0] _334;
    wire [7:0] _335;
    wire [15:0] _336;
    wire [31:0] _338;
    wire [16:0] _330;
    wire [2:0] _327;
    wire [6:0] _328;
    wire _323;
    wire [1:0] _324;
    wire [3:0] _325;
    wire [7:0] _326;
    wire [14:0] _329;
    wire [31:0] _331;
    wire [17:0] _321;
    wire [5:0] _319;
    wire _315;
    wire [1:0] _316;
    wire [3:0] _317;
    wire [7:0] _318;
    wire [13:0] _320;
    wire [31:0] _322;
    wire [18:0] _313;
    wire [4:0] _311;
    wire _307;
    wire [1:0] _308;
    wire [3:0] _309;
    wire [7:0] _310;
    wire [12:0] _312;
    wire [31:0] _314;
    wire [19:0] _305;
    wire _300;
    wire [1:0] _301;
    wire [3:0] _302;
    wire [7:0] _303;
    wire [11:0] _304;
    wire [31:0] _306;
    wire [20:0] _298;
    wire [2:0] _296;
    wire _292;
    wire [1:0] _293;
    wire [3:0] _294;
    wire [7:0] _295;
    wire [10:0] _297;
    wire [31:0] _299;
    wire [21:0] _290;
    wire _285;
    wire [1:0] _286;
    wire [3:0] _287;
    wire [7:0] _288;
    wire [9:0] _289;
    wire [31:0] _291;
    wire [22:0] _283;
    wire _278;
    wire [1:0] _279;
    wire [3:0] _280;
    wire [7:0] _281;
    wire [8:0] _282;
    wire [31:0] _284;
    wire [23:0] _276;
    wire _272;
    wire [1:0] _273;
    wire [3:0] _274;
    wire [7:0] _275;
    wire [31:0] _277;
    wire [24:0] _270;
    wire [2:0] _268;
    wire _265;
    wire [1:0] _266;
    wire [3:0] _267;
    wire [6:0] _269;
    wire [31:0] _271;
    wire [25:0] _263;
    wire _259;
    wire [1:0] _260;
    wire [3:0] _261;
    wire [5:0] _262;
    wire [31:0] _264;
    wire [26:0] _257;
    wire _253;
    wire [1:0] _254;
    wire [3:0] _255;
    wire [4:0] _256;
    wire [31:0] _258;
    wire [27:0] _251;
    wire _248;
    wire [1:0] _249;
    wire [3:0] _250;
    wire [31:0] _252;
    wire [28:0] _246;
    wire _243;
    wire [1:0] _244;
    wire [2:0] _245;
    wire [31:0] _247;
    wire [29:0] _241;
    wire _239;
    wire [1:0] _240;
    wire [31:0] _242;
    wire [30:0] _237;
    wire _236;
    wire [31:0] _238;
    reg [31:0] _476;
    wire [31:0] _234 = 32'b00000000000000000000000000011111;
    wire _235;
    wire [31:0] _478;
    wire [31:0] _232 = 32'b00000000000000000000000000000000;
    wire _229;
    wire [30:0] _228 = 31'b0000000000000000000000000000000;
    wire [31:0] _230;
    wire [1:0] _226;
    wire [29:0] _225 = 30'b000000000000000000000000000000;
    wire [31:0] _227;
    wire [2:0] _223;
    wire [28:0] _222 = 29'b00000000000000000000000000000;
    wire [31:0] _224;
    wire [3:0] _220;
    wire [27:0] _219 = 28'b0000000000000000000000000000;
    wire [31:0] _221;
    wire [4:0] _217;
    wire [26:0] _216 = 27'b000000000000000000000000000;
    wire [31:0] _218;
    wire [5:0] _214;
    wire [25:0] _213 = 26'b00000000000000000000000000;
    wire [31:0] _215;
    wire [6:0] _211;
    wire [24:0] _210 = 25'b0000000000000000000000000;
    wire [31:0] _212;
    wire [7:0] _208;
    wire [23:0] _207 = 24'b000000000000000000000000;
    wire [31:0] _209;
    wire [8:0] _205;
    wire [22:0] _204 = 23'b00000000000000000000000;
    wire [31:0] _206;
    wire [9:0] _202;
    wire [21:0] _201 = 22'b0000000000000000000000;
    wire [31:0] _203;
    wire [10:0] _199;
    wire [20:0] _198 = 21'b000000000000000000000;
    wire [31:0] _200;
    wire [11:0] _196;
    wire [19:0] _195 = 20'b00000000000000000000;
    wire [31:0] _197;
    wire [12:0] _193;
    wire [18:0] _192 = 19'b0000000000000000000;
    wire [31:0] _194;
    wire [13:0] _190;
    wire [17:0] _189 = 18'b000000000000000000;
    wire [31:0] _191;
    wire [14:0] _187;
    wire [16:0] _186 = 17'b00000000000000000;
    wire [31:0] _188;
    wire [15:0] _184;
    wire [15:0] _183 = 16'b0000000000000000;
    wire [31:0] _185;
    wire [16:0] _181;
    wire [14:0] _180 = 15'b000000000000000;
    wire [31:0] _182;
    wire [17:0] _178;
    wire [13:0] _177 = 14'b00000000000000;
    wire [31:0] _179;
    wire [18:0] _175;
    wire [12:0] _174 = 13'b0000000000000;
    wire [31:0] _176;
    wire [19:0] _172;
    wire [11:0] _171 = 12'b000000000000;
    wire [31:0] _173;
    wire [20:0] _169;
    wire [10:0] _168 = 11'b00000000000;
    wire [31:0] _170;
    wire [21:0] _166;
    wire [9:0] _165 = 10'b0000000000;
    wire [31:0] _167;
    wire [22:0] _163;
    wire [8:0] _162 = 9'b000000000;
    wire [31:0] _164;
    wire [23:0] _160;
    wire [7:0] _159 = 8'b00000000;
    wire [31:0] _161;
    wire [24:0] _157;
    wire [6:0] _156 = 7'b0000000;
    wire [31:0] _158;
    wire [25:0] _154;
    wire [5:0] _153 = 6'b000000;
    wire [31:0] _155;
    wire [26:0] _151;
    wire [4:0] _150 = 5'b00000;
    wire [31:0] _152;
    wire [27:0] _148;
    wire [3:0] _147 = 4'b0000;
    wire [31:0] _149;
    wire [28:0] _145;
    wire [2:0] _144 = 3'b000;
    wire [31:0] _146;
    wire [29:0] _142;
    wire [1:0] _141 = 2'b00;
    wire [31:0] _143;
    wire [30:0] _139;
    wire _138 = 1'b0;
    wire [31:0] _140;
    reg [31:0] _231;
    wire [31:0] _136 = 32'b00000000000000000000000000011111;
    wire _137;
    wire [31:0] _233;
    wire [6:0] _3;
    wire _135;
    wire [31:0] _479;
    wire [31:0] _134;
    wire _132;
    wire [30:0] _131 = 31'b0000000000000000000000000000000;
    wire [31:0] _133;
    wire [30:0] _127;
    wire _125;
    wire _126;
    wire [31:0] _128;
    wire [30:0] _123;
    wire _121;
    wire _122;
    wire [31:0] _124;
    wire _129;
    wire [30:0] _120 = 31'b0000000000000000000000000000000;
    wire [31:0] _130;
    wire [31:0] _118 = 32'b00000000000000000000000000000000;
    wire [30:0] _115 = 31'b0000000000000000000000000000000;
    wire _114;
    wire [31:0] _116;
    wire [29:0] _112 = 30'b000000000000000000000000000000;
    wire [1:0] _111;
    wire [31:0] _113;
    wire [28:0] _109 = 29'b00000000000000000000000000000;
    wire [2:0] _108;
    wire [31:0] _110;
    wire [27:0] _106 = 28'b0000000000000000000000000000;
    wire [3:0] _105;
    wire [31:0] _107;
    wire [26:0] _103 = 27'b000000000000000000000000000;
    wire [4:0] _102;
    wire [31:0] _104;
    wire [25:0] _100 = 26'b00000000000000000000000000;
    wire [5:0] _99;
    wire [31:0] _101;
    wire [24:0] _97 = 25'b0000000000000000000000000;
    wire [6:0] _96;
    wire [31:0] _98;
    wire [23:0] _94 = 24'b000000000000000000000000;
    wire [7:0] _93;
    wire [31:0] _95;
    wire [22:0] _91 = 23'b00000000000000000000000;
    wire [8:0] _90;
    wire [31:0] _92;
    wire [21:0] _88 = 22'b0000000000000000000000;
    wire [9:0] _87;
    wire [31:0] _89;
    wire [20:0] _85 = 21'b000000000000000000000;
    wire [10:0] _84;
    wire [31:0] _86;
    wire [19:0] _82 = 20'b00000000000000000000;
    wire [11:0] _81;
    wire [31:0] _83;
    wire [18:0] _79 = 19'b0000000000000000000;
    wire [12:0] _78;
    wire [31:0] _80;
    wire [17:0] _76 = 18'b000000000000000000;
    wire [13:0] _75;
    wire [31:0] _77;
    wire [16:0] _73 = 17'b00000000000000000;
    wire [14:0] _72;
    wire [31:0] _74;
    wire [15:0] _70 = 16'b0000000000000000;
    wire [15:0] _69;
    wire [31:0] _71;
    wire [14:0] _67 = 15'b000000000000000;
    wire [16:0] _66;
    wire [31:0] _68;
    wire [13:0] _64 = 14'b00000000000000;
    wire [17:0] _63;
    wire [31:0] _65;
    wire [12:0] _61 = 13'b0000000000000;
    wire [18:0] _60;
    wire [31:0] _62;
    wire [11:0] _58 = 12'b000000000000;
    wire [19:0] _57;
    wire [31:0] _59;
    wire [10:0] _55 = 11'b00000000000;
    wire [20:0] _54;
    wire [31:0] _56;
    wire [9:0] _52 = 10'b0000000000;
    wire [21:0] _51;
    wire [31:0] _53;
    wire [8:0] _49 = 9'b000000000;
    wire [22:0] _48;
    wire [31:0] _50;
    wire [7:0] _46 = 8'b00000000;
    wire [23:0] _45;
    wire [31:0] _47;
    wire [6:0] _43 = 7'b0000000;
    wire [24:0] _42;
    wire [31:0] _44;
    wire [5:0] _40 = 6'b000000;
    wire [25:0] _39;
    wire [31:0] _41;
    wire [4:0] _37 = 5'b00000;
    wire [26:0] _36;
    wire [31:0] _38;
    wire [3:0] _34 = 4'b0000;
    wire [27:0] _33;
    wire [31:0] _35;
    wire [2:0] _31 = 3'b000;
    wire [28:0] _30;
    wire [31:0] _32;
    wire [1:0] _28 = 2'b00;
    wire [29:0] _27;
    wire [31:0] _29;
    wire _25 = 1'b0;
    wire [30:0] _24;
    wire [31:0] _26;
    reg [31:0] _117;
    wire [31:0] _22 = 32'b00000000000000000000000000011111;
    wire _23;
    wire [31:0] _119;
    wire [31:0] _5;
    wire [31:0] _7;
    wire [31:0] _21;
    wire [2:0] _9;
    reg [31:0] _482;

    /* logic */
    assign _17 = _16 < _3;
    always @* begin
        case (_9)
        0: _20 <= _11;
        1: _20 <= _12;
        2: _20 <= _13;
        3: _20 <= _14;
        4: _20 <= _15;
        5: _20 <= _17;
        6: _20 <= _18;
        default: _20 <= _19;
        endcase
    end
    assign _481 = _7 & _5;
    assign _480 = _7 | _5;
    assign _474 = _7[31:31];
    assign _470 = { _466, _465 };
    assign _471 = { _467, _470 };
    assign _472 = { _468, _471 };
    assign _465 = _7[31:31];
    assign _466 = { _465, _465 };
    assign _467 = { _466, _466 };
    assign _468 = { _467, _467 };
    assign _469 = { _468, _468 };
    assign _473 = { _469, _472 };
    assign _475 = { _473, _474 };
    assign _463 = _7[31:30];
    assign _460 = { _457, _456 };
    assign _461 = { _458, _460 };
    assign _455 = _7[31:31];
    assign _456 = { _455, _455 };
    assign _457 = { _456, _456 };
    assign _458 = { _457, _457 };
    assign _459 = { _458, _458 };
    assign _462 = { _459, _461 };
    assign _464 = { _462, _463 };
    assign _453 = _7[31:29];
    assign _450 = { _447, _445 };
    assign _451 = { _448, _450 };
    assign _445 = _7[31:31];
    assign _446 = { _445, _445 };
    assign _447 = { _446, _446 };
    assign _448 = { _447, _447 };
    assign _449 = { _448, _448 };
    assign _452 = { _449, _451 };
    assign _454 = { _452, _453 };
    assign _443 = _7[31:28];
    assign _441 = { _439, _438 };
    assign _436 = _7[31:31];
    assign _437 = { _436, _436 };
    assign _438 = { _437, _437 };
    assign _439 = { _438, _438 };
    assign _440 = { _439, _439 };
    assign _442 = { _440, _441 };
    assign _444 = { _442, _443 };
    assign _434 = _7[31:27];
    assign _431 = { _427, _426 };
    assign _432 = { _429, _431 };
    assign _426 = _7[31:31];
    assign _427 = { _426, _426 };
    assign _428 = { _427, _427 };
    assign _429 = { _428, _428 };
    assign _430 = { _429, _429 };
    assign _433 = { _430, _432 };
    assign _435 = { _433, _434 };
    assign _424 = _7[31:26];
    assign _422 = { _420, _418 };
    assign _417 = _7[31:31];
    assign _418 = { _417, _417 };
    assign _419 = { _418, _418 };
    assign _420 = { _419, _419 };
    assign _421 = { _420, _420 };
    assign _423 = { _421, _422 };
    assign _425 = { _423, _424 };
    assign _415 = _7[31:25];
    assign _413 = { _411, _408 };
    assign _408 = _7[31:31];
    assign _409 = { _408, _408 };
    assign _410 = { _409, _409 };
    assign _411 = { _410, _410 };
    assign _412 = { _411, _411 };
    assign _414 = { _412, _413 };
    assign _416 = { _414, _415 };
    assign _406 = _7[31:24];
    assign _400 = _7[31:31];
    assign _401 = { _400, _400 };
    assign _402 = { _401, _401 };
    assign _403 = { _402, _402 };
    assign _404 = { _403, _403 };
    assign _405 = { _404, _403 };
    assign _407 = { _405, _406 };
    assign _398 = _7[31:23];
    assign _395 = { _391, _390 };
    assign _396 = { _392, _395 };
    assign _390 = _7[31:31];
    assign _391 = { _390, _390 };
    assign _392 = { _391, _391 };
    assign _393 = { _392, _392 };
    assign _394 = { _393, _393 };
    assign _397 = { _394, _396 };
    assign _399 = { _397, _398 };
    assign _388 = _7[31:22];
    assign _386 = { _383, _382 };
    assign _381 = _7[31:31];
    assign _382 = { _381, _381 };
    assign _383 = { _382, _382 };
    assign _384 = { _383, _383 };
    assign _385 = { _384, _384 };
    assign _387 = { _385, _386 };
    assign _389 = { _387, _388 };
    assign _379 = _7[31:21];
    assign _377 = { _374, _372 };
    assign _372 = _7[31:31];
    assign _373 = { _372, _372 };
    assign _374 = { _373, _373 };
    assign _375 = { _374, _374 };
    assign _376 = { _375, _375 };
    assign _378 = { _376, _377 };
    assign _380 = { _378, _379 };
    assign _370 = _7[31:20];
    assign _364 = _7[31:31];
    assign _365 = { _364, _364 };
    assign _366 = { _365, _365 };
    assign _367 = { _366, _366 };
    assign _368 = { _367, _367 };
    assign _369 = { _368, _366 };
    assign _371 = { _369, _370 };
    assign _362 = _7[31:19];
    assign _360 = { _356, _355 };
    assign _355 = _7[31:31];
    assign _356 = { _355, _355 };
    assign _357 = { _356, _356 };
    assign _358 = { _357, _357 };
    assign _359 = { _358, _358 };
    assign _361 = { _359, _360 };
    assign _363 = { _361, _362 };
    assign _353 = _7[31:18];
    assign _347 = _7[31:31];
    assign _348 = { _347, _347 };
    assign _349 = { _348, _348 };
    assign _350 = { _349, _349 };
    assign _351 = { _350, _350 };
    assign _352 = { _351, _348 };
    assign _354 = { _352, _353 };
    assign _345 = _7[31:17];
    assign _339 = _7[31:31];
    assign _340 = { _339, _339 };
    assign _341 = { _340, _340 };
    assign _342 = { _341, _341 };
    assign _343 = { _342, _342 };
    assign _344 = { _343, _339 };
    assign _346 = { _344, _345 };
    assign _337 = _7[31:16];
    assign _332 = _7[31:31];
    assign _333 = { _332, _332 };
    assign _334 = { _333, _333 };
    assign _335 = { _334, _334 };
    assign _336 = { _335, _335 };
    assign _338 = { _336, _337 };
    assign _330 = _7[31:15];
    assign _327 = { _324, _323 };
    assign _328 = { _325, _327 };
    assign _323 = _7[31:31];
    assign _324 = { _323, _323 };
    assign _325 = { _324, _324 };
    assign _326 = { _325, _325 };
    assign _329 = { _326, _328 };
    assign _331 = { _329, _330 };
    assign _321 = _7[31:14];
    assign _319 = { _317, _316 };
    assign _315 = _7[31:31];
    assign _316 = { _315, _315 };
    assign _317 = { _316, _316 };
    assign _318 = { _317, _317 };
    assign _320 = { _318, _319 };
    assign _322 = { _320, _321 };
    assign _313 = _7[31:13];
    assign _311 = { _309, _307 };
    assign _307 = _7[31:31];
    assign _308 = { _307, _307 };
    assign _309 = { _308, _308 };
    assign _310 = { _309, _309 };
    assign _312 = { _310, _311 };
    assign _314 = { _312, _313 };
    assign _305 = _7[31:12];
    assign _300 = _7[31:31];
    assign _301 = { _300, _300 };
    assign _302 = { _301, _301 };
    assign _303 = { _302, _302 };
    assign _304 = { _303, _302 };
    assign _306 = { _304, _305 };
    assign _298 = _7[31:11];
    assign _296 = { _293, _292 };
    assign _292 = _7[31:31];
    assign _293 = { _292, _292 };
    assign _294 = { _293, _293 };
    assign _295 = { _294, _294 };
    assign _297 = { _295, _296 };
    assign _299 = { _297, _298 };
    assign _290 = _7[31:10];
    assign _285 = _7[31:31];
    assign _286 = { _285, _285 };
    assign _287 = { _286, _286 };
    assign _288 = { _287, _287 };
    assign _289 = { _288, _286 };
    assign _291 = { _289, _290 };
    assign _283 = _7[31:9];
    assign _278 = _7[31:31];
    assign _279 = { _278, _278 };
    assign _280 = { _279, _279 };
    assign _281 = { _280, _280 };
    assign _282 = { _281, _278 };
    assign _284 = { _282, _283 };
    assign _276 = _7[31:8];
    assign _272 = _7[31:31];
    assign _273 = { _272, _272 };
    assign _274 = { _273, _273 };
    assign _275 = { _274, _274 };
    assign _277 = { _275, _276 };
    assign _270 = _7[31:7];
    assign _268 = { _266, _265 };
    assign _265 = _7[31:31];
    assign _266 = { _265, _265 };
    assign _267 = { _266, _266 };
    assign _269 = { _267, _268 };
    assign _271 = { _269, _270 };
    assign _263 = _7[31:6];
    assign _259 = _7[31:31];
    assign _260 = { _259, _259 };
    assign _261 = { _260, _260 };
    assign _262 = { _261, _260 };
    assign _264 = { _262, _263 };
    assign _257 = _7[31:5];
    assign _253 = _7[31:31];
    assign _254 = { _253, _253 };
    assign _255 = { _254, _254 };
    assign _256 = { _255, _253 };
    assign _258 = { _256, _257 };
    assign _251 = _7[31:4];
    assign _248 = _7[31:31];
    assign _249 = { _248, _248 };
    assign _250 = { _249, _249 };
    assign _252 = { _250, _251 };
    assign _246 = _7[31:3];
    assign _243 = _7[31:31];
    assign _244 = { _243, _243 };
    assign _245 = { _244, _243 };
    assign _247 = { _245, _246 };
    assign _241 = _7[31:2];
    assign _239 = _7[31:31];
    assign _240 = { _239, _239 };
    assign _242 = { _240, _241 };
    assign _237 = _7[31:1];
    assign _236 = _7[31:31];
    assign _238 = { _236, _237 };
    always @* begin
        case (_5)
        0: _476 <= _7;
        1: _476 <= _238;
        2: _476 <= _242;
        3: _476 <= _247;
        4: _476 <= _252;
        5: _476 <= _258;
        6: _476 <= _264;
        7: _476 <= _271;
        8: _476 <= _277;
        9: _476 <= _284;
        10: _476 <= _291;
        11: _476 <= _299;
        12: _476 <= _306;
        13: _476 <= _314;
        14: _476 <= _322;
        15: _476 <= _331;
        16: _476 <= _338;
        17: _476 <= _346;
        18: _476 <= _354;
        19: _476 <= _363;
        20: _476 <= _371;
        21: _476 <= _380;
        22: _476 <= _389;
        23: _476 <= _399;
        24: _476 <= _407;
        25: _476 <= _416;
        26: _476 <= _425;
        27: _476 <= _435;
        28: _476 <= _444;
        29: _476 <= _454;
        30: _476 <= _464;
        default: _476 <= _475;
        endcase
    end
    assign _235 = _234 < _5;
    assign _478 = _235 ? _477 : _476;
    assign _229 = _7[31:31];
    assign _230 = { _228, _229 };
    assign _226 = _7[31:30];
    assign _227 = { _225, _226 };
    assign _223 = _7[31:29];
    assign _224 = { _222, _223 };
    assign _220 = _7[31:28];
    assign _221 = { _219, _220 };
    assign _217 = _7[31:27];
    assign _218 = { _216, _217 };
    assign _214 = _7[31:26];
    assign _215 = { _213, _214 };
    assign _211 = _7[31:25];
    assign _212 = { _210, _211 };
    assign _208 = _7[31:24];
    assign _209 = { _207, _208 };
    assign _205 = _7[31:23];
    assign _206 = { _204, _205 };
    assign _202 = _7[31:22];
    assign _203 = { _201, _202 };
    assign _199 = _7[31:21];
    assign _200 = { _198, _199 };
    assign _196 = _7[31:20];
    assign _197 = { _195, _196 };
    assign _193 = _7[31:19];
    assign _194 = { _192, _193 };
    assign _190 = _7[31:18];
    assign _191 = { _189, _190 };
    assign _187 = _7[31:17];
    assign _188 = { _186, _187 };
    assign _184 = _7[31:16];
    assign _185 = { _183, _184 };
    assign _181 = _7[31:15];
    assign _182 = { _180, _181 };
    assign _178 = _7[31:14];
    assign _179 = { _177, _178 };
    assign _175 = _7[31:13];
    assign _176 = { _174, _175 };
    assign _172 = _7[31:12];
    assign _173 = { _171, _172 };
    assign _169 = _7[31:11];
    assign _170 = { _168, _169 };
    assign _166 = _7[31:10];
    assign _167 = { _165, _166 };
    assign _163 = _7[31:9];
    assign _164 = { _162, _163 };
    assign _160 = _7[31:8];
    assign _161 = { _159, _160 };
    assign _157 = _7[31:7];
    assign _158 = { _156, _157 };
    assign _154 = _7[31:6];
    assign _155 = { _153, _154 };
    assign _151 = _7[31:5];
    assign _152 = { _150, _151 };
    assign _148 = _7[31:4];
    assign _149 = { _147, _148 };
    assign _145 = _7[31:3];
    assign _146 = { _144, _145 };
    assign _142 = _7[31:2];
    assign _143 = { _141, _142 };
    assign _139 = _7[31:1];
    assign _140 = { _138, _139 };
    always @* begin
        case (_5)
        0: _231 <= _7;
        1: _231 <= _140;
        2: _231 <= _143;
        3: _231 <= _146;
        4: _231 <= _149;
        5: _231 <= _152;
        6: _231 <= _155;
        7: _231 <= _158;
        8: _231 <= _161;
        9: _231 <= _164;
        10: _231 <= _167;
        11: _231 <= _170;
        12: _231 <= _173;
        13: _231 <= _176;
        14: _231 <= _179;
        15: _231 <= _182;
        16: _231 <= _185;
        17: _231 <= _188;
        18: _231 <= _191;
        19: _231 <= _194;
        20: _231 <= _197;
        21: _231 <= _200;
        22: _231 <= _203;
        23: _231 <= _206;
        24: _231 <= _209;
        25: _231 <= _212;
        26: _231 <= _215;
        27: _231 <= _218;
        28: _231 <= _221;
        29: _231 <= _224;
        30: _231 <= _227;
        default: _231 <= _230;
        endcase
    end
    assign _137 = _136 < _5;
    assign _233 = _137 ? _232 : _231;
    assign _3 = funct7;
    assign _135 = _3[0:0];
    assign _479 = _135 ? _478 : _233;
    assign _134 = _7 ^ _5;
    assign _132 = _7 < _5;
    assign _133 = { _131, _132 };
    assign _127 = _5[30:0];
    assign _125 = _5[31:31];
    assign _126 = ~ _125;
    assign _128 = { _126, _127 };
    assign _123 = _7[30:0];
    assign _121 = _7[31:31];
    assign _122 = ~ _121;
    assign _124 = { _122, _123 };
    assign _129 = _124 < _128;
    assign _130 = { _120, _129 };
    assign _114 = _7[0:0];
    assign _116 = { _114, _115 };
    assign _111 = _7[1:0];
    assign _113 = { _111, _112 };
    assign _108 = _7[2:0];
    assign _110 = { _108, _109 };
    assign _105 = _7[3:0];
    assign _107 = { _105, _106 };
    assign _102 = _7[4:0];
    assign _104 = { _102, _103 };
    assign _99 = _7[5:0];
    assign _101 = { _99, _100 };
    assign _96 = _7[6:0];
    assign _98 = { _96, _97 };
    assign _93 = _7[7:0];
    assign _95 = { _93, _94 };
    assign _90 = _7[8:0];
    assign _92 = { _90, _91 };
    assign _87 = _7[9:0];
    assign _89 = { _87, _88 };
    assign _84 = _7[10:0];
    assign _86 = { _84, _85 };
    assign _81 = _7[11:0];
    assign _83 = { _81, _82 };
    assign _78 = _7[12:0];
    assign _80 = { _78, _79 };
    assign _75 = _7[13:0];
    assign _77 = { _75, _76 };
    assign _72 = _7[14:0];
    assign _74 = { _72, _73 };
    assign _69 = _7[15:0];
    assign _71 = { _69, _70 };
    assign _66 = _7[16:0];
    assign _68 = { _66, _67 };
    assign _63 = _7[17:0];
    assign _65 = { _63, _64 };
    assign _60 = _7[18:0];
    assign _62 = { _60, _61 };
    assign _57 = _7[19:0];
    assign _59 = { _57, _58 };
    assign _54 = _7[20:0];
    assign _56 = { _54, _55 };
    assign _51 = _7[21:0];
    assign _53 = { _51, _52 };
    assign _48 = _7[22:0];
    assign _50 = { _48, _49 };
    assign _45 = _7[23:0];
    assign _47 = { _45, _46 };
    assign _42 = _7[24:0];
    assign _44 = { _42, _43 };
    assign _39 = _7[25:0];
    assign _41 = { _39, _40 };
    assign _36 = _7[26:0];
    assign _38 = { _36, _37 };
    assign _33 = _7[27:0];
    assign _35 = { _33, _34 };
    assign _30 = _7[28:0];
    assign _32 = { _30, _31 };
    assign _27 = _7[29:0];
    assign _29 = { _27, _28 };
    assign _24 = _7[30:0];
    assign _26 = { _24, _25 };
    always @* begin
        case (_5)
        0: _117 <= _7;
        1: _117 <= _26;
        2: _117 <= _29;
        3: _117 <= _32;
        4: _117 <= _35;
        5: _117 <= _38;
        6: _117 <= _41;
        7: _117 <= _44;
        8: _117 <= _47;
        9: _117 <= _50;
        10: _117 <= _53;
        11: _117 <= _56;
        12: _117 <= _59;
        13: _117 <= _62;
        14: _117 <= _65;
        15: _117 <= _68;
        16: _117 <= _71;
        17: _117 <= _74;
        18: _117 <= _77;
        19: _117 <= _80;
        20: _117 <= _83;
        21: _117 <= _86;
        22: _117 <= _89;
        23: _117 <= _92;
        24: _117 <= _95;
        25: _117 <= _98;
        26: _117 <= _101;
        27: _117 <= _104;
        28: _117 <= _107;
        29: _117 <= _110;
        30: _117 <= _113;
        default: _117 <= _116;
        endcase
    end
    assign _23 = _22 < _5;
    assign _119 = _23 ? _118 : _117;
    assign _5 = rhs;
    assign _7 = lhs;
    assign _21 = _7 + _5;
    assign _9 = funct3;
    always @* begin
        case (_9)
        0: _482 <= _21;
        1: _482 <= _119;
        2: _482 <= _130;
        3: _482 <= _133;
        4: _482 <= _134;
        5: _482 <= _479;
        6: _482 <= _480;
        default: _482 <= _481;
        endcase
    end

    /* aliases */

    /* output assignments */
    assign new_rd = _482;
    assign error = _20;

endmodule
