module Uart_tx (
    uart_rx,
    clear,
    clock,
    data_out_valid,
    data_out,
    parity_error,
    stop_bit_unstable
);

    input uart_rx;
    input clear;
    input clock;
    output data_out_valid;
    output [7:0] data_out;
    output parity_error;
    output stop_bit_unstable;

    /* signal declarations */
    wire _48;
    wire _49;
    wire _50;
    wire _30 = 1'b0;
    wire _29;
    wire _51;
    wire _2;
    wire [7:0] _57 = 8'b00000000;
    wire [7:0] _56 = 8'b00000000;
    wire [7:0] _177 = 8'b00000000;
    wire _172;
    wire _171;
    wire _170;
    wire _169;
    wire _168;
    wire _167;
    wire [6:0] _160;
    wire [5:0] _161;
    wire [4:0] _162;
    wire [3:0] _163;
    wire [2:0] _164;
    wire [1:0] _165;
    wire _166;
    wire [7:0] _173;
    wire _158;
    wire _157;
    wire _156;
    wire _155;
    wire _154;
    wire _153;
    wire [6:0] _146;
    wire [5:0] _147;
    wire [4:0] _148;
    wire [3:0] _149;
    wire [2:0] _150;
    wire [1:0] _151;
    wire _152;
    wire [7:0] _159;
    wire _144;
    wire _143;
    wire _142;
    wire _141;
    wire _140;
    wire _139;
    wire [6:0] _132;
    wire [5:0] _133;
    wire [4:0] _134;
    wire [3:0] _135;
    wire [2:0] _136;
    wire [1:0] _137;
    wire _138;
    wire [7:0] _145;
    wire _130;
    wire _129;
    wire _128;
    wire _127;
    wire _126;
    wire _125;
    wire [6:0] _118;
    wire [5:0] _119;
    wire [4:0] _120;
    wire [3:0] _121;
    wire [2:0] _122;
    wire [1:0] _123;
    wire _124;
    wire [7:0] _131;
    wire _116;
    wire _115;
    wire _114;
    wire _113;
    wire _112;
    wire _111;
    wire [6:0] _104;
    wire [5:0] _105;
    wire [4:0] _106;
    wire [3:0] _107;
    wire [2:0] _108;
    wire [1:0] _109;
    wire _110;
    wire [7:0] _117;
    wire _102;
    wire _101;
    wire _100;
    wire _99;
    wire _98;
    wire _97;
    wire [6:0] _90;
    wire [5:0] _91;
    wire [4:0] _92;
    wire [3:0] _93;
    wire [2:0] _94;
    wire [1:0] _95;
    wire _96;
    wire [7:0] _103;
    wire _88;
    wire _87;
    wire _86;
    wire _85;
    wire _84;
    wire _83;
    wire [6:0] _76;
    wire [5:0] _77;
    wire [4:0] _78;
    wire [3:0] _79;
    wire [2:0] _80;
    wire [1:0] _81;
    wire _82;
    wire [7:0] _89;
    wire _74;
    wire _73;
    wire _72;
    wire _71;
    wire _70;
    wire _69;
    wire [6:0] _62;
    wire [5:0] _63;
    wire [4:0] _64;
    wire [3:0] _65;
    wire [2:0] _66;
    wire [1:0] _67;
    wire _68;
    wire [7:0] _75;
    reg [7:0] data_with_new_bit;
    wire [7:0] _175;
    wire _55;
    wire [7:0] _176;
    wire _53;
    wire [7:0] _178;
    wire [7:0] _4;
    reg [7:0] _58;
    wire _45 = 1'b0;
    wire _44 = 1'b0;
    wire _184 = 1'b0;
    wire _182;
    wire _181;
    wire _183;
    wire _179;
    wire _185;
    wire _6;
    reg rx_parity_bit;
    wire _42 = 1'b0;
    wire _41 = 1'b0;
    wire _191 = 1'b0;
    wire _188;
    wire _189;
    wire _187;
    wire _190;
    wire _186;
    wire _192;
    wire _7;
    reg calculated_parity_bit;
    wire _47;
    wire _22 = 1'b0;
    wire _21 = 1'b0;
    wire _201 = 1'b0;
    wire _197 = 1'b1;
    wire _195 = 1'b0;
    wire _196;
    wire _198;
    wire _199;
    wire _194;
    wire _200;
    wire _193;
    wire _202;
    wire _8;
    reg _24;
    wire _246;
    wire _247;
    wire _248;
    wire _249;
    wire _245 = 1'b0;
    wire [1:0] _26 = 2'b00;
    wire [1:0] _25 = 2'b00;
    wire _239 = 1'b0;
    wire _10;
    wire _240;
    wire _241;
    wire [1:0] _242;
    wire [2:0] _234 = 3'b111;
    wire [2:0] _60 = 3'b000;
    wire [2:0] _59 = 3'b000;
    wire [2:0] _209 = 3'b000;
    wire [2:0] _205 = 3'b001;
    wire [2:0] _206;
    wire [2:0] _207;
    wire _204;
    wire [2:0] _208;
    wire _203;
    wire [2:0] _210;
    wire [2:0] _11;
    reg [2:0] which_data_bit;
    wire _235;
    wire [1:0] _236;
    wire [1:0] _237;
    wire [1:0] _232;
    wire [1:0] _39 = 2'b01;
    wire [1:0] _37 = 2'b00;
    wire [1:0] _36 = 2'b00;
    wire [1:0] _217 = 2'b00;
    wire [1:0] _213 = 2'b01;
    wire [1:0] _214;
    wire [1:0] _215;
    wire _212;
    wire [1:0] _216;
    wire _211;
    wire [1:0] _218;
    wire [1:0] _12;
    reg [1:0] _38;
    wire _40;
    wire [1:0] _229;
    wire [4:0] _34 = 5'b00000;
    wire vdd = 1'b1;
    wire [4:0] _32 = 5'b00000;
    wire _14;
    wire [4:0] _31 = 5'b00000;
    wire _16;
    wire [4:0] _223 = 5'b00000;
    wire [4:0] _221 = 5'b00001;
    wire [4:0] _222;
    wire [4:0] _219 = 5'b10001;
    wire _220;
    wire [4:0] _224;
    wire [4:0] _17;
    reg [4:0] _33;
    wire switch_cycle;
    wire [1:0] _230;
    wire [1:0] _28 = 2'b11;
    wire _228;
    wire [1:0] _231;
    wire [1:0] _180 = 2'b10;
    wire _227;
    wire [1:0] _233;
    wire [1:0] _54 = 2'b01;
    wire _226;
    wire [1:0] _238;
    wire [1:0] _52 = 2'b00;
    wire _225;
    wire [1:0] _243;
    wire [1:0] _18;
    reg [1:0] current_state;
    wire _244;
    wire _250;
    wire _19;

    /* logic */
    assign _48 = ~ _47;
    assign _49 = _40 ? _48 : _30;
    assign _50 = switch_cycle ? _49 : _30;
    assign _29 = current_state == _28;
    assign _51 = _29 ? _50 : _30;
    assign _2 = _51;
    assign _172 = _58[0:0];
    assign _171 = _160[0:0];
    assign _170 = _161[0:0];
    assign _169 = _162[0:0];
    assign _168 = _163[0:0];
    assign _167 = _164[0:0];
    assign _160 = _58[7:1];
    assign _161 = _160[6:1];
    assign _162 = _161[5:1];
    assign _163 = _162[4:1];
    assign _164 = _163[3:1];
    assign _165 = _164[2:1];
    assign _166 = _165[0:0];
    assign _173 = { _10, _166, _167, _168, _169, _170, _171, _172 };
    assign _158 = _58[0:0];
    assign _157 = _146[0:0];
    assign _156 = _147[0:0];
    assign _155 = _148[0:0];
    assign _154 = _149[0:0];
    assign _153 = _150[0:0];
    assign _146 = _58[7:1];
    assign _147 = _146[6:1];
    assign _148 = _147[5:1];
    assign _149 = _148[4:1];
    assign _150 = _149[3:1];
    assign _151 = _150[2:1];
    assign _152 = _151[1:1];
    assign _159 = { _152, _10, _153, _154, _155, _156, _157, _158 };
    assign _144 = _58[0:0];
    assign _143 = _132[0:0];
    assign _142 = _133[0:0];
    assign _141 = _134[0:0];
    assign _140 = _135[0:0];
    assign _139 = _137[0:0];
    assign _132 = _58[7:1];
    assign _133 = _132[6:1];
    assign _134 = _133[5:1];
    assign _135 = _134[4:1];
    assign _136 = _135[3:1];
    assign _137 = _136[2:1];
    assign _138 = _137[1:1];
    assign _145 = { _138, _139, _10, _140, _141, _142, _143, _144 };
    assign _130 = _58[0:0];
    assign _129 = _118[0:0];
    assign _128 = _119[0:0];
    assign _127 = _120[0:0];
    assign _126 = _122[0:0];
    assign _125 = _123[0:0];
    assign _118 = _58[7:1];
    assign _119 = _118[6:1];
    assign _120 = _119[5:1];
    assign _121 = _120[4:1];
    assign _122 = _121[3:1];
    assign _123 = _122[2:1];
    assign _124 = _123[1:1];
    assign _131 = { _124, _125, _126, _10, _127, _128, _129, _130 };
    assign _116 = _58[0:0];
    assign _115 = _104[0:0];
    assign _114 = _105[0:0];
    assign _113 = _107[0:0];
    assign _112 = _108[0:0];
    assign _111 = _109[0:0];
    assign _104 = _58[7:1];
    assign _105 = _104[6:1];
    assign _106 = _105[5:1];
    assign _107 = _106[4:1];
    assign _108 = _107[3:1];
    assign _109 = _108[2:1];
    assign _110 = _109[1:1];
    assign _117 = { _110, _111, _112, _113, _10, _114, _115, _116 };
    assign _102 = _58[0:0];
    assign _101 = _90[0:0];
    assign _100 = _92[0:0];
    assign _99 = _93[0:0];
    assign _98 = _94[0:0];
    assign _97 = _95[0:0];
    assign _90 = _58[7:1];
    assign _91 = _90[6:1];
    assign _92 = _91[5:1];
    assign _93 = _92[4:1];
    assign _94 = _93[3:1];
    assign _95 = _94[2:1];
    assign _96 = _95[1:1];
    assign _103 = { _96, _97, _98, _99, _100, _10, _101, _102 };
    assign _88 = _58[0:0];
    assign _87 = _77[0:0];
    assign _86 = _78[0:0];
    assign _85 = _79[0:0];
    assign _84 = _80[0:0];
    assign _83 = _81[0:0];
    assign _76 = _58[7:1];
    assign _77 = _76[6:1];
    assign _78 = _77[5:1];
    assign _79 = _78[4:1];
    assign _80 = _79[3:1];
    assign _81 = _80[2:1];
    assign _82 = _81[1:1];
    assign _89 = { _82, _83, _84, _85, _86, _87, _10, _88 };
    assign _74 = _62[0:0];
    assign _73 = _63[0:0];
    assign _72 = _64[0:0];
    assign _71 = _65[0:0];
    assign _70 = _66[0:0];
    assign _69 = _67[0:0];
    assign _62 = _58[7:1];
    assign _63 = _62[6:1];
    assign _64 = _63[5:1];
    assign _65 = _64[4:1];
    assign _66 = _65[3:1];
    assign _67 = _66[2:1];
    assign _68 = _67[1:1];
    assign _75 = { _68, _69, _70, _71, _72, _73, _74, _10 };
    always @* begin
        case (which_data_bit)
        0: data_with_new_bit <= _75;
        1: data_with_new_bit <= _89;
        2: data_with_new_bit <= _103;
        3: data_with_new_bit <= _117;
        4: data_with_new_bit <= _131;
        5: data_with_new_bit <= _145;
        6: data_with_new_bit <= _159;
        default: data_with_new_bit <= _173;
        endcase
    end
    assign _175 = switch_cycle ? data_with_new_bit : _58;
    assign _55 = current_state == _54;
    assign _176 = _55 ? _175 : _58;
    assign _53 = current_state == _52;
    assign _178 = _53 ? _177 : _176;
    assign _4 = _178;
    always @(posedge _16) begin
        _58 <= _4;
    end
    assign _182 = switch_cycle ? _10 : rx_parity_bit;
    assign _181 = current_state == _180;
    assign _183 = _181 ? _182 : rx_parity_bit;
    assign _179 = current_state == _52;
    assign _185 = _179 ? _184 : _183;
    assign _6 = _185;
    always @(posedge _16) begin
        rx_parity_bit <= _6;
    end
    assign _188 = calculated_parity_bit + _10;
    assign _189 = switch_cycle ? _188 : calculated_parity_bit;
    assign _187 = current_state == _54;
    assign _190 = _187 ? _189 : calculated_parity_bit;
    assign _186 = current_state == _52;
    assign _192 = _186 ? _191 : _190;
    assign _7 = _192;
    always @(posedge _16) begin
        calculated_parity_bit <= _7;
    end
    assign _47 = calculated_parity_bit == rx_parity_bit;
    assign _196 = _10 == _195;
    assign _198 = _196 ? _197 : _24;
    assign _199 = switch_cycle ? _198 : _24;
    assign _194 = current_state == _28;
    assign _200 = _194 ? _199 : _24;
    assign _193 = current_state == _52;
    assign _202 = _193 ? _201 : _200;
    assign _8 = _202;
    always @(posedge _16) begin
        _24 <= _8;
    end
    assign _246 = ~ _24;
    assign _247 = _246 & _47;
    assign _248 = _40 ? _247 : _245;
    assign _249 = switch_cycle ? _248 : _245;
    assign _10 = uart_rx;
    assign _240 = _10 == _239;
    assign _241 = switch_cycle & _240;
    assign _242 = _241 ? _54 : current_state;
    assign _206 = which_data_bit + _205;
    assign _207 = switch_cycle ? _206 : which_data_bit;
    assign _204 = current_state == _54;
    assign _208 = _204 ? _207 : which_data_bit;
    assign _203 = current_state == _52;
    assign _210 = _203 ? _209 : _208;
    assign _11 = _210;
    always @(posedge _16) begin
        which_data_bit <= _11;
    end
    assign _235 = which_data_bit == _234;
    assign _236 = _235 ? _180 : current_state;
    assign _237 = switch_cycle ? _236 : current_state;
    assign _232 = switch_cycle ? _28 : current_state;
    assign _214 = _38 + _213;
    assign _215 = switch_cycle ? _214 : _38;
    assign _212 = current_state == _28;
    assign _216 = _212 ? _215 : _38;
    assign _211 = current_state == _52;
    assign _218 = _211 ? _217 : _216;
    assign _12 = _218;
    always @(posedge _16) begin
        _38 <= _12;
    end
    assign _40 = _38 == _39;
    assign _229 = _40 ? _52 : current_state;
    assign _14 = clear;
    assign _16 = clock;
    assign _222 = _33 + _221;
    assign _220 = _33 == _219;
    assign _224 = _220 ? _223 : _222;
    assign _17 = _224;
    always @(posedge _16) begin
        if (_14)
            _33 <= _32;
        else
            _33 <= _17;
    end
    assign switch_cycle = _33 == _34;
    assign _230 = switch_cycle ? _229 : current_state;
    assign _228 = current_state == _28;
    assign _231 = _228 ? _230 : current_state;
    assign _227 = current_state == _180;
    assign _233 = _227 ? _232 : _231;
    assign _226 = current_state == _54;
    assign _238 = _226 ? _237 : _233;
    assign _225 = current_state == _52;
    assign _243 = _225 ? _242 : _238;
    assign _18 = _243;
    always @(posedge _16) begin
        if (_14)
            current_state <= _26;
        else
            current_state <= _18;
    end
    assign _244 = current_state == _28;
    assign _250 = _244 ? _249 : _245;
    assign _19 = _250;

    /* aliases */

    /* output assignments */
    assign data_out_valid = _19;
    assign data_out = _58;
    assign parity_error = _2;
    assign stop_bit_unstable = _24;

endmodule
