module Op_0 (
    rhs,
    lhs,
    funct7,
    funct3,
    new_rd,
    error
);

    input [31:0] rhs;
    input [31:0] lhs;
    input [6:0] funct7;
    input [2:0] funct3;
    output [31:0] new_rd;
    output error;

    /* signal declarations */
    wire _20 = 1'b0;
    wire _19 = 1'b0;
    wire [6:0] _17 = 7'b0000001;
    wire _18;
    wire _16 = 1'b0;
    wire _15 = 1'b0;
    wire _14 = 1'b0;
    wire _13 = 1'b0;
    wire [6:0] _11 = 7'b0000001;
    wire _12;
    reg _21;
    wire [31:0] _485;
    wire [31:0] _484;
    wire [31:0] _481 = 32'b11111111111111111111111111111111;
    wire _478;
    wire [2:0] _474;
    wire [6:0] _475;
    wire [14:0] _476;
    wire _469;
    wire [1:0] _470;
    wire [3:0] _471;
    wire [7:0] _472;
    wire [15:0] _473;
    wire [30:0] _477;
    wire [31:0] _479;
    wire [1:0] _467;
    wire [5:0] _464;
    wire [13:0] _465;
    wire _459;
    wire [1:0] _460;
    wire [3:0] _461;
    wire [7:0] _462;
    wire [15:0] _463;
    wire [29:0] _466;
    wire [31:0] _468;
    wire [2:0] _457;
    wire [4:0] _454;
    wire [12:0] _455;
    wire _449;
    wire [1:0] _450;
    wire [3:0] _451;
    wire [7:0] _452;
    wire [15:0] _453;
    wire [28:0] _456;
    wire [31:0] _458;
    wire [3:0] _447;
    wire [11:0] _445;
    wire _440;
    wire [1:0] _441;
    wire [3:0] _442;
    wire [7:0] _443;
    wire [15:0] _444;
    wire [27:0] _446;
    wire [31:0] _448;
    wire [4:0] _438;
    wire [2:0] _435;
    wire [10:0] _436;
    wire _430;
    wire [1:0] _431;
    wire [3:0] _432;
    wire [7:0] _433;
    wire [15:0] _434;
    wire [26:0] _437;
    wire [31:0] _439;
    wire [5:0] _428;
    wire [9:0] _426;
    wire _421;
    wire [1:0] _422;
    wire [3:0] _423;
    wire [7:0] _424;
    wire [15:0] _425;
    wire [25:0] _427;
    wire [31:0] _429;
    wire [6:0] _419;
    wire [8:0] _417;
    wire _412;
    wire [1:0] _413;
    wire [3:0] _414;
    wire [7:0] _415;
    wire [15:0] _416;
    wire [24:0] _418;
    wire [31:0] _420;
    wire [7:0] _410;
    wire _404;
    wire [1:0] _405;
    wire [3:0] _406;
    wire [7:0] _407;
    wire [15:0] _408;
    wire [23:0] _409;
    wire [31:0] _411;
    wire [8:0] _402;
    wire [2:0] _399;
    wire [6:0] _400;
    wire _394;
    wire [1:0] _395;
    wire [3:0] _396;
    wire [7:0] _397;
    wire [15:0] _398;
    wire [22:0] _401;
    wire [31:0] _403;
    wire [9:0] _392;
    wire [5:0] _390;
    wire _385;
    wire [1:0] _386;
    wire [3:0] _387;
    wire [7:0] _388;
    wire [15:0] _389;
    wire [21:0] _391;
    wire [31:0] _393;
    wire [10:0] _383;
    wire [4:0] _381;
    wire _376;
    wire [1:0] _377;
    wire [3:0] _378;
    wire [7:0] _379;
    wire [15:0] _380;
    wire [20:0] _382;
    wire [31:0] _384;
    wire [11:0] _374;
    wire _368;
    wire [1:0] _369;
    wire [3:0] _370;
    wire [7:0] _371;
    wire [15:0] _372;
    wire [19:0] _373;
    wire [31:0] _375;
    wire [12:0] _366;
    wire [2:0] _364;
    wire _359;
    wire [1:0] _360;
    wire [3:0] _361;
    wire [7:0] _362;
    wire [15:0] _363;
    wire [18:0] _365;
    wire [31:0] _367;
    wire [13:0] _357;
    wire _351;
    wire [1:0] _352;
    wire [3:0] _353;
    wire [7:0] _354;
    wire [15:0] _355;
    wire [17:0] _356;
    wire [31:0] _358;
    wire [14:0] _349;
    wire _343;
    wire [1:0] _344;
    wire [3:0] _345;
    wire [7:0] _346;
    wire [15:0] _347;
    wire [16:0] _348;
    wire [31:0] _350;
    wire [15:0] _341;
    wire _336;
    wire [1:0] _337;
    wire [3:0] _338;
    wire [7:0] _339;
    wire [15:0] _340;
    wire [31:0] _342;
    wire [16:0] _334;
    wire [2:0] _331;
    wire [6:0] _332;
    wire _327;
    wire [1:0] _328;
    wire [3:0] _329;
    wire [7:0] _330;
    wire [14:0] _333;
    wire [31:0] _335;
    wire [17:0] _325;
    wire [5:0] _323;
    wire _319;
    wire [1:0] _320;
    wire [3:0] _321;
    wire [7:0] _322;
    wire [13:0] _324;
    wire [31:0] _326;
    wire [18:0] _317;
    wire [4:0] _315;
    wire _311;
    wire [1:0] _312;
    wire [3:0] _313;
    wire [7:0] _314;
    wire [12:0] _316;
    wire [31:0] _318;
    wire [19:0] _309;
    wire _304;
    wire [1:0] _305;
    wire [3:0] _306;
    wire [7:0] _307;
    wire [11:0] _308;
    wire [31:0] _310;
    wire [20:0] _302;
    wire [2:0] _300;
    wire _296;
    wire [1:0] _297;
    wire [3:0] _298;
    wire [7:0] _299;
    wire [10:0] _301;
    wire [31:0] _303;
    wire [21:0] _294;
    wire _289;
    wire [1:0] _290;
    wire [3:0] _291;
    wire [7:0] _292;
    wire [9:0] _293;
    wire [31:0] _295;
    wire [22:0] _287;
    wire _282;
    wire [1:0] _283;
    wire [3:0] _284;
    wire [7:0] _285;
    wire [8:0] _286;
    wire [31:0] _288;
    wire [23:0] _280;
    wire _276;
    wire [1:0] _277;
    wire [3:0] _278;
    wire [7:0] _279;
    wire [31:0] _281;
    wire [24:0] _274;
    wire [2:0] _272;
    wire _269;
    wire [1:0] _270;
    wire [3:0] _271;
    wire [6:0] _273;
    wire [31:0] _275;
    wire [25:0] _267;
    wire _263;
    wire [1:0] _264;
    wire [3:0] _265;
    wire [5:0] _266;
    wire [31:0] _268;
    wire [26:0] _261;
    wire _257;
    wire [1:0] _258;
    wire [3:0] _259;
    wire [4:0] _260;
    wire [31:0] _262;
    wire [27:0] _255;
    wire _252;
    wire [1:0] _253;
    wire [3:0] _254;
    wire [31:0] _256;
    wire [28:0] _250;
    wire _247;
    wire [1:0] _248;
    wire [2:0] _249;
    wire [31:0] _251;
    wire [29:0] _245;
    wire _243;
    wire [1:0] _244;
    wire [31:0] _246;
    wire [30:0] _241;
    wire _240;
    wire [31:0] _242;
    reg [31:0] _480;
    wire [31:0] _238 = 32'b00000000000000000000000000011111;
    wire _239;
    wire [31:0] _482;
    wire [31:0] _236 = 32'b00000000000000000000000000000000;
    wire _233;
    wire [30:0] _232 = 31'b0000000000000000000000000000000;
    wire [31:0] _234;
    wire [1:0] _230;
    wire [29:0] _229 = 30'b000000000000000000000000000000;
    wire [31:0] _231;
    wire [2:0] _227;
    wire [28:0] _226 = 29'b00000000000000000000000000000;
    wire [31:0] _228;
    wire [3:0] _224;
    wire [27:0] _223 = 28'b0000000000000000000000000000;
    wire [31:0] _225;
    wire [4:0] _221;
    wire [26:0] _220 = 27'b000000000000000000000000000;
    wire [31:0] _222;
    wire [5:0] _218;
    wire [25:0] _217 = 26'b00000000000000000000000000;
    wire [31:0] _219;
    wire [6:0] _215;
    wire [24:0] _214 = 25'b0000000000000000000000000;
    wire [31:0] _216;
    wire [7:0] _212;
    wire [23:0] _211 = 24'b000000000000000000000000;
    wire [31:0] _213;
    wire [8:0] _209;
    wire [22:0] _208 = 23'b00000000000000000000000;
    wire [31:0] _210;
    wire [9:0] _206;
    wire [21:0] _205 = 22'b0000000000000000000000;
    wire [31:0] _207;
    wire [10:0] _203;
    wire [20:0] _202 = 21'b000000000000000000000;
    wire [31:0] _204;
    wire [11:0] _200;
    wire [19:0] _199 = 20'b00000000000000000000;
    wire [31:0] _201;
    wire [12:0] _197;
    wire [18:0] _196 = 19'b0000000000000000000;
    wire [31:0] _198;
    wire [13:0] _194;
    wire [17:0] _193 = 18'b000000000000000000;
    wire [31:0] _195;
    wire [14:0] _191;
    wire [16:0] _190 = 17'b00000000000000000;
    wire [31:0] _192;
    wire [15:0] _188;
    wire [15:0] _187 = 16'b0000000000000000;
    wire [31:0] _189;
    wire [16:0] _185;
    wire [14:0] _184 = 15'b000000000000000;
    wire [31:0] _186;
    wire [17:0] _182;
    wire [13:0] _181 = 14'b00000000000000;
    wire [31:0] _183;
    wire [18:0] _179;
    wire [12:0] _178 = 13'b0000000000000;
    wire [31:0] _180;
    wire [19:0] _176;
    wire [11:0] _175 = 12'b000000000000;
    wire [31:0] _177;
    wire [20:0] _173;
    wire [10:0] _172 = 11'b00000000000;
    wire [31:0] _174;
    wire [21:0] _170;
    wire [9:0] _169 = 10'b0000000000;
    wire [31:0] _171;
    wire [22:0] _167;
    wire [8:0] _166 = 9'b000000000;
    wire [31:0] _168;
    wire [23:0] _164;
    wire [7:0] _163 = 8'b00000000;
    wire [31:0] _165;
    wire [24:0] _161;
    wire [6:0] _160 = 7'b0000000;
    wire [31:0] _162;
    wire [25:0] _158;
    wire [5:0] _157 = 6'b000000;
    wire [31:0] _159;
    wire [26:0] _155;
    wire [4:0] _154 = 5'b00000;
    wire [31:0] _156;
    wire [27:0] _152;
    wire [3:0] _151 = 4'b0000;
    wire [31:0] _153;
    wire [28:0] _149;
    wire [2:0] _148 = 3'b000;
    wire [31:0] _150;
    wire [29:0] _146;
    wire [1:0] _145 = 2'b00;
    wire [31:0] _147;
    wire [30:0] _143;
    wire _142 = 1'b0;
    wire [31:0] _144;
    reg [31:0] _235;
    wire [31:0] _140 = 32'b00000000000000000000000000011111;
    wire _141;
    wire [31:0] _237;
    wire _139;
    wire [31:0] _483;
    wire [31:0] _138;
    wire _136;
    wire [30:0] _135 = 31'b0000000000000000000000000000000;
    wire [31:0] _137;
    wire [30:0] _131;
    wire _129;
    wire _130;
    wire [31:0] _132;
    wire [30:0] _127;
    wire _125;
    wire _126;
    wire [31:0] _128;
    wire _133;
    wire [30:0] _124 = 31'b0000000000000000000000000000000;
    wire [31:0] _134;
    wire [31:0] _122 = 32'b00000000000000000000000000000000;
    wire [30:0] _119 = 31'b0000000000000000000000000000000;
    wire _118;
    wire [31:0] _120;
    wire [29:0] _116 = 30'b000000000000000000000000000000;
    wire [1:0] _115;
    wire [31:0] _117;
    wire [28:0] _113 = 29'b00000000000000000000000000000;
    wire [2:0] _112;
    wire [31:0] _114;
    wire [27:0] _110 = 28'b0000000000000000000000000000;
    wire [3:0] _109;
    wire [31:0] _111;
    wire [26:0] _107 = 27'b000000000000000000000000000;
    wire [4:0] _106;
    wire [31:0] _108;
    wire [25:0] _104 = 26'b00000000000000000000000000;
    wire [5:0] _103;
    wire [31:0] _105;
    wire [24:0] _101 = 25'b0000000000000000000000000;
    wire [6:0] _100;
    wire [31:0] _102;
    wire [23:0] _98 = 24'b000000000000000000000000;
    wire [7:0] _97;
    wire [31:0] _99;
    wire [22:0] _95 = 23'b00000000000000000000000;
    wire [8:0] _94;
    wire [31:0] _96;
    wire [21:0] _92 = 22'b0000000000000000000000;
    wire [9:0] _91;
    wire [31:0] _93;
    wire [20:0] _89 = 21'b000000000000000000000;
    wire [10:0] _88;
    wire [31:0] _90;
    wire [19:0] _86 = 20'b00000000000000000000;
    wire [11:0] _85;
    wire [31:0] _87;
    wire [18:0] _83 = 19'b0000000000000000000;
    wire [12:0] _82;
    wire [31:0] _84;
    wire [17:0] _80 = 18'b000000000000000000;
    wire [13:0] _79;
    wire [31:0] _81;
    wire [16:0] _77 = 17'b00000000000000000;
    wire [14:0] _76;
    wire [31:0] _78;
    wire [15:0] _74 = 16'b0000000000000000;
    wire [15:0] _73;
    wire [31:0] _75;
    wire [14:0] _71 = 15'b000000000000000;
    wire [16:0] _70;
    wire [31:0] _72;
    wire [13:0] _68 = 14'b00000000000000;
    wire [17:0] _67;
    wire [31:0] _69;
    wire [12:0] _65 = 13'b0000000000000;
    wire [18:0] _64;
    wire [31:0] _66;
    wire [11:0] _62 = 12'b000000000000;
    wire [19:0] _61;
    wire [31:0] _63;
    wire [10:0] _59 = 11'b00000000000;
    wire [20:0] _58;
    wire [31:0] _60;
    wire [9:0] _56 = 10'b0000000000;
    wire [21:0] _55;
    wire [31:0] _57;
    wire [8:0] _53 = 9'b000000000;
    wire [22:0] _52;
    wire [31:0] _54;
    wire [7:0] _50 = 8'b00000000;
    wire [23:0] _49;
    wire [31:0] _51;
    wire [6:0] _47 = 7'b0000000;
    wire [24:0] _46;
    wire [31:0] _48;
    wire [5:0] _44 = 6'b000000;
    wire [25:0] _43;
    wire [31:0] _45;
    wire [4:0] _41 = 5'b00000;
    wire [26:0] _40;
    wire [31:0] _42;
    wire [3:0] _38 = 4'b0000;
    wire [27:0] _37;
    wire [31:0] _39;
    wire [2:0] _35 = 3'b000;
    wire [28:0] _34;
    wire [31:0] _36;
    wire [1:0] _32 = 2'b00;
    wire [29:0] _31;
    wire [31:0] _33;
    wire _29 = 1'b0;
    wire [30:0] _28;
    wire [31:0] _30;
    reg [31:0] _121;
    wire [31:0] _26 = 32'b00000000000000000000000000011111;
    wire _27;
    wire [31:0] _123;
    wire [31:0] _24;
    wire [31:0] _3;
    wire [31:0] _5;
    wire [31:0] _23;
    wire [6:0] _7;
    wire _22;
    wire [31:0] _25;
    wire [2:0] _9;
    reg [31:0] _486;

    /* logic */
    assign _18 = _17 < _7;
    assign _12 = _11 < _7;
    always @* begin
        case (_9)
        0: _21 <= _12;
        1: _21 <= _13;
        2: _21 <= _14;
        3: _21 <= _15;
        4: _21 <= _16;
        5: _21 <= _18;
        6: _21 <= _19;
        default: _21 <= _20;
        endcase
    end
    assign _485 = _5 & _3;
    assign _484 = _5 | _3;
    assign _478 = _5[31:31];
    assign _474 = { _470, _469 };
    assign _475 = { _471, _474 };
    assign _476 = { _472, _475 };
    assign _469 = _5[31:31];
    assign _470 = { _469, _469 };
    assign _471 = { _470, _470 };
    assign _472 = { _471, _471 };
    assign _473 = { _472, _472 };
    assign _477 = { _473, _476 };
    assign _479 = { _477, _478 };
    assign _467 = _5[31:30];
    assign _464 = { _461, _460 };
    assign _465 = { _462, _464 };
    assign _459 = _5[31:31];
    assign _460 = { _459, _459 };
    assign _461 = { _460, _460 };
    assign _462 = { _461, _461 };
    assign _463 = { _462, _462 };
    assign _466 = { _463, _465 };
    assign _468 = { _466, _467 };
    assign _457 = _5[31:29];
    assign _454 = { _451, _449 };
    assign _455 = { _452, _454 };
    assign _449 = _5[31:31];
    assign _450 = { _449, _449 };
    assign _451 = { _450, _450 };
    assign _452 = { _451, _451 };
    assign _453 = { _452, _452 };
    assign _456 = { _453, _455 };
    assign _458 = { _456, _457 };
    assign _447 = _5[31:28];
    assign _445 = { _443, _442 };
    assign _440 = _5[31:31];
    assign _441 = { _440, _440 };
    assign _442 = { _441, _441 };
    assign _443 = { _442, _442 };
    assign _444 = { _443, _443 };
    assign _446 = { _444, _445 };
    assign _448 = { _446, _447 };
    assign _438 = _5[31:27];
    assign _435 = { _431, _430 };
    assign _436 = { _433, _435 };
    assign _430 = _5[31:31];
    assign _431 = { _430, _430 };
    assign _432 = { _431, _431 };
    assign _433 = { _432, _432 };
    assign _434 = { _433, _433 };
    assign _437 = { _434, _436 };
    assign _439 = { _437, _438 };
    assign _428 = _5[31:26];
    assign _426 = { _424, _422 };
    assign _421 = _5[31:31];
    assign _422 = { _421, _421 };
    assign _423 = { _422, _422 };
    assign _424 = { _423, _423 };
    assign _425 = { _424, _424 };
    assign _427 = { _425, _426 };
    assign _429 = { _427, _428 };
    assign _419 = _5[31:25];
    assign _417 = { _415, _412 };
    assign _412 = _5[31:31];
    assign _413 = { _412, _412 };
    assign _414 = { _413, _413 };
    assign _415 = { _414, _414 };
    assign _416 = { _415, _415 };
    assign _418 = { _416, _417 };
    assign _420 = { _418, _419 };
    assign _410 = _5[31:24];
    assign _404 = _5[31:31];
    assign _405 = { _404, _404 };
    assign _406 = { _405, _405 };
    assign _407 = { _406, _406 };
    assign _408 = { _407, _407 };
    assign _409 = { _408, _407 };
    assign _411 = { _409, _410 };
    assign _402 = _5[31:23];
    assign _399 = { _395, _394 };
    assign _400 = { _396, _399 };
    assign _394 = _5[31:31];
    assign _395 = { _394, _394 };
    assign _396 = { _395, _395 };
    assign _397 = { _396, _396 };
    assign _398 = { _397, _397 };
    assign _401 = { _398, _400 };
    assign _403 = { _401, _402 };
    assign _392 = _5[31:22];
    assign _390 = { _387, _386 };
    assign _385 = _5[31:31];
    assign _386 = { _385, _385 };
    assign _387 = { _386, _386 };
    assign _388 = { _387, _387 };
    assign _389 = { _388, _388 };
    assign _391 = { _389, _390 };
    assign _393 = { _391, _392 };
    assign _383 = _5[31:21];
    assign _381 = { _378, _376 };
    assign _376 = _5[31:31];
    assign _377 = { _376, _376 };
    assign _378 = { _377, _377 };
    assign _379 = { _378, _378 };
    assign _380 = { _379, _379 };
    assign _382 = { _380, _381 };
    assign _384 = { _382, _383 };
    assign _374 = _5[31:20];
    assign _368 = _5[31:31];
    assign _369 = { _368, _368 };
    assign _370 = { _369, _369 };
    assign _371 = { _370, _370 };
    assign _372 = { _371, _371 };
    assign _373 = { _372, _370 };
    assign _375 = { _373, _374 };
    assign _366 = _5[31:19];
    assign _364 = { _360, _359 };
    assign _359 = _5[31:31];
    assign _360 = { _359, _359 };
    assign _361 = { _360, _360 };
    assign _362 = { _361, _361 };
    assign _363 = { _362, _362 };
    assign _365 = { _363, _364 };
    assign _367 = { _365, _366 };
    assign _357 = _5[31:18];
    assign _351 = _5[31:31];
    assign _352 = { _351, _351 };
    assign _353 = { _352, _352 };
    assign _354 = { _353, _353 };
    assign _355 = { _354, _354 };
    assign _356 = { _355, _352 };
    assign _358 = { _356, _357 };
    assign _349 = _5[31:17];
    assign _343 = _5[31:31];
    assign _344 = { _343, _343 };
    assign _345 = { _344, _344 };
    assign _346 = { _345, _345 };
    assign _347 = { _346, _346 };
    assign _348 = { _347, _343 };
    assign _350 = { _348, _349 };
    assign _341 = _5[31:16];
    assign _336 = _5[31:31];
    assign _337 = { _336, _336 };
    assign _338 = { _337, _337 };
    assign _339 = { _338, _338 };
    assign _340 = { _339, _339 };
    assign _342 = { _340, _341 };
    assign _334 = _5[31:15];
    assign _331 = { _328, _327 };
    assign _332 = { _329, _331 };
    assign _327 = _5[31:31];
    assign _328 = { _327, _327 };
    assign _329 = { _328, _328 };
    assign _330 = { _329, _329 };
    assign _333 = { _330, _332 };
    assign _335 = { _333, _334 };
    assign _325 = _5[31:14];
    assign _323 = { _321, _320 };
    assign _319 = _5[31:31];
    assign _320 = { _319, _319 };
    assign _321 = { _320, _320 };
    assign _322 = { _321, _321 };
    assign _324 = { _322, _323 };
    assign _326 = { _324, _325 };
    assign _317 = _5[31:13];
    assign _315 = { _313, _311 };
    assign _311 = _5[31:31];
    assign _312 = { _311, _311 };
    assign _313 = { _312, _312 };
    assign _314 = { _313, _313 };
    assign _316 = { _314, _315 };
    assign _318 = { _316, _317 };
    assign _309 = _5[31:12];
    assign _304 = _5[31:31];
    assign _305 = { _304, _304 };
    assign _306 = { _305, _305 };
    assign _307 = { _306, _306 };
    assign _308 = { _307, _306 };
    assign _310 = { _308, _309 };
    assign _302 = _5[31:11];
    assign _300 = { _297, _296 };
    assign _296 = _5[31:31];
    assign _297 = { _296, _296 };
    assign _298 = { _297, _297 };
    assign _299 = { _298, _298 };
    assign _301 = { _299, _300 };
    assign _303 = { _301, _302 };
    assign _294 = _5[31:10];
    assign _289 = _5[31:31];
    assign _290 = { _289, _289 };
    assign _291 = { _290, _290 };
    assign _292 = { _291, _291 };
    assign _293 = { _292, _290 };
    assign _295 = { _293, _294 };
    assign _287 = _5[31:9];
    assign _282 = _5[31:31];
    assign _283 = { _282, _282 };
    assign _284 = { _283, _283 };
    assign _285 = { _284, _284 };
    assign _286 = { _285, _282 };
    assign _288 = { _286, _287 };
    assign _280 = _5[31:8];
    assign _276 = _5[31:31];
    assign _277 = { _276, _276 };
    assign _278 = { _277, _277 };
    assign _279 = { _278, _278 };
    assign _281 = { _279, _280 };
    assign _274 = _5[31:7];
    assign _272 = { _270, _269 };
    assign _269 = _5[31:31];
    assign _270 = { _269, _269 };
    assign _271 = { _270, _270 };
    assign _273 = { _271, _272 };
    assign _275 = { _273, _274 };
    assign _267 = _5[31:6];
    assign _263 = _5[31:31];
    assign _264 = { _263, _263 };
    assign _265 = { _264, _264 };
    assign _266 = { _265, _264 };
    assign _268 = { _266, _267 };
    assign _261 = _5[31:5];
    assign _257 = _5[31:31];
    assign _258 = { _257, _257 };
    assign _259 = { _258, _258 };
    assign _260 = { _259, _257 };
    assign _262 = { _260, _261 };
    assign _255 = _5[31:4];
    assign _252 = _5[31:31];
    assign _253 = { _252, _252 };
    assign _254 = { _253, _253 };
    assign _256 = { _254, _255 };
    assign _250 = _5[31:3];
    assign _247 = _5[31:31];
    assign _248 = { _247, _247 };
    assign _249 = { _248, _247 };
    assign _251 = { _249, _250 };
    assign _245 = _5[31:2];
    assign _243 = _5[31:31];
    assign _244 = { _243, _243 };
    assign _246 = { _244, _245 };
    assign _241 = _5[31:1];
    assign _240 = _5[31:31];
    assign _242 = { _240, _241 };
    always @* begin
        case (_3)
        0: _480 <= _5;
        1: _480 <= _242;
        2: _480 <= _246;
        3: _480 <= _251;
        4: _480 <= _256;
        5: _480 <= _262;
        6: _480 <= _268;
        7: _480 <= _275;
        8: _480 <= _281;
        9: _480 <= _288;
        10: _480 <= _295;
        11: _480 <= _303;
        12: _480 <= _310;
        13: _480 <= _318;
        14: _480 <= _326;
        15: _480 <= _335;
        16: _480 <= _342;
        17: _480 <= _350;
        18: _480 <= _358;
        19: _480 <= _367;
        20: _480 <= _375;
        21: _480 <= _384;
        22: _480 <= _393;
        23: _480 <= _403;
        24: _480 <= _411;
        25: _480 <= _420;
        26: _480 <= _429;
        27: _480 <= _439;
        28: _480 <= _448;
        29: _480 <= _458;
        30: _480 <= _468;
        default: _480 <= _479;
        endcase
    end
    assign _239 = _238 < _3;
    assign _482 = _239 ? _481 : _480;
    assign _233 = _5[31:31];
    assign _234 = { _232, _233 };
    assign _230 = _5[31:30];
    assign _231 = { _229, _230 };
    assign _227 = _5[31:29];
    assign _228 = { _226, _227 };
    assign _224 = _5[31:28];
    assign _225 = { _223, _224 };
    assign _221 = _5[31:27];
    assign _222 = { _220, _221 };
    assign _218 = _5[31:26];
    assign _219 = { _217, _218 };
    assign _215 = _5[31:25];
    assign _216 = { _214, _215 };
    assign _212 = _5[31:24];
    assign _213 = { _211, _212 };
    assign _209 = _5[31:23];
    assign _210 = { _208, _209 };
    assign _206 = _5[31:22];
    assign _207 = { _205, _206 };
    assign _203 = _5[31:21];
    assign _204 = { _202, _203 };
    assign _200 = _5[31:20];
    assign _201 = { _199, _200 };
    assign _197 = _5[31:19];
    assign _198 = { _196, _197 };
    assign _194 = _5[31:18];
    assign _195 = { _193, _194 };
    assign _191 = _5[31:17];
    assign _192 = { _190, _191 };
    assign _188 = _5[31:16];
    assign _189 = { _187, _188 };
    assign _185 = _5[31:15];
    assign _186 = { _184, _185 };
    assign _182 = _5[31:14];
    assign _183 = { _181, _182 };
    assign _179 = _5[31:13];
    assign _180 = { _178, _179 };
    assign _176 = _5[31:12];
    assign _177 = { _175, _176 };
    assign _173 = _5[31:11];
    assign _174 = { _172, _173 };
    assign _170 = _5[31:10];
    assign _171 = { _169, _170 };
    assign _167 = _5[31:9];
    assign _168 = { _166, _167 };
    assign _164 = _5[31:8];
    assign _165 = { _163, _164 };
    assign _161 = _5[31:7];
    assign _162 = { _160, _161 };
    assign _158 = _5[31:6];
    assign _159 = { _157, _158 };
    assign _155 = _5[31:5];
    assign _156 = { _154, _155 };
    assign _152 = _5[31:4];
    assign _153 = { _151, _152 };
    assign _149 = _5[31:3];
    assign _150 = { _148, _149 };
    assign _146 = _5[31:2];
    assign _147 = { _145, _146 };
    assign _143 = _5[31:1];
    assign _144 = { _142, _143 };
    always @* begin
        case (_3)
        0: _235 <= _5;
        1: _235 <= _144;
        2: _235 <= _147;
        3: _235 <= _150;
        4: _235 <= _153;
        5: _235 <= _156;
        6: _235 <= _159;
        7: _235 <= _162;
        8: _235 <= _165;
        9: _235 <= _168;
        10: _235 <= _171;
        11: _235 <= _174;
        12: _235 <= _177;
        13: _235 <= _180;
        14: _235 <= _183;
        15: _235 <= _186;
        16: _235 <= _189;
        17: _235 <= _192;
        18: _235 <= _195;
        19: _235 <= _198;
        20: _235 <= _201;
        21: _235 <= _204;
        22: _235 <= _207;
        23: _235 <= _210;
        24: _235 <= _213;
        25: _235 <= _216;
        26: _235 <= _219;
        27: _235 <= _222;
        28: _235 <= _225;
        29: _235 <= _228;
        30: _235 <= _231;
        default: _235 <= _234;
        endcase
    end
    assign _141 = _140 < _3;
    assign _237 = _141 ? _236 : _235;
    assign _139 = _7[0:0];
    assign _483 = _139 ? _482 : _237;
    assign _138 = _5 ^ _3;
    assign _136 = _5 < _3;
    assign _137 = { _135, _136 };
    assign _131 = _3[30:0];
    assign _129 = _3[31:31];
    assign _130 = ~ _129;
    assign _132 = { _130, _131 };
    assign _127 = _5[30:0];
    assign _125 = _5[31:31];
    assign _126 = ~ _125;
    assign _128 = { _126, _127 };
    assign _133 = _128 < _132;
    assign _134 = { _124, _133 };
    assign _118 = _5[0:0];
    assign _120 = { _118, _119 };
    assign _115 = _5[1:0];
    assign _117 = { _115, _116 };
    assign _112 = _5[2:0];
    assign _114 = { _112, _113 };
    assign _109 = _5[3:0];
    assign _111 = { _109, _110 };
    assign _106 = _5[4:0];
    assign _108 = { _106, _107 };
    assign _103 = _5[5:0];
    assign _105 = { _103, _104 };
    assign _100 = _5[6:0];
    assign _102 = { _100, _101 };
    assign _97 = _5[7:0];
    assign _99 = { _97, _98 };
    assign _94 = _5[8:0];
    assign _96 = { _94, _95 };
    assign _91 = _5[9:0];
    assign _93 = { _91, _92 };
    assign _88 = _5[10:0];
    assign _90 = { _88, _89 };
    assign _85 = _5[11:0];
    assign _87 = { _85, _86 };
    assign _82 = _5[12:0];
    assign _84 = { _82, _83 };
    assign _79 = _5[13:0];
    assign _81 = { _79, _80 };
    assign _76 = _5[14:0];
    assign _78 = { _76, _77 };
    assign _73 = _5[15:0];
    assign _75 = { _73, _74 };
    assign _70 = _5[16:0];
    assign _72 = { _70, _71 };
    assign _67 = _5[17:0];
    assign _69 = { _67, _68 };
    assign _64 = _5[18:0];
    assign _66 = { _64, _65 };
    assign _61 = _5[19:0];
    assign _63 = { _61, _62 };
    assign _58 = _5[20:0];
    assign _60 = { _58, _59 };
    assign _55 = _5[21:0];
    assign _57 = { _55, _56 };
    assign _52 = _5[22:0];
    assign _54 = { _52, _53 };
    assign _49 = _5[23:0];
    assign _51 = { _49, _50 };
    assign _46 = _5[24:0];
    assign _48 = { _46, _47 };
    assign _43 = _5[25:0];
    assign _45 = { _43, _44 };
    assign _40 = _5[26:0];
    assign _42 = { _40, _41 };
    assign _37 = _5[27:0];
    assign _39 = { _37, _38 };
    assign _34 = _5[28:0];
    assign _36 = { _34, _35 };
    assign _31 = _5[29:0];
    assign _33 = { _31, _32 };
    assign _28 = _5[30:0];
    assign _30 = { _28, _29 };
    always @* begin
        case (_3)
        0: _121 <= _5;
        1: _121 <= _30;
        2: _121 <= _33;
        3: _121 <= _36;
        4: _121 <= _39;
        5: _121 <= _42;
        6: _121 <= _45;
        7: _121 <= _48;
        8: _121 <= _51;
        9: _121 <= _54;
        10: _121 <= _57;
        11: _121 <= _60;
        12: _121 <= _63;
        13: _121 <= _66;
        14: _121 <= _69;
        15: _121 <= _72;
        16: _121 <= _75;
        17: _121 <= _78;
        18: _121 <= _81;
        19: _121 <= _84;
        20: _121 <= _87;
        21: _121 <= _90;
        22: _121 <= _93;
        23: _121 <= _96;
        24: _121 <= _99;
        25: _121 <= _102;
        26: _121 <= _105;
        27: _121 <= _108;
        28: _121 <= _111;
        29: _121 <= _114;
        30: _121 <= _117;
        default: _121 <= _120;
        endcase
    end
    assign _27 = _26 < _3;
    assign _123 = _27 ? _122 : _121;
    assign _24 = _5 + _3;
    assign _3 = rhs;
    assign _5 = lhs;
    assign _23 = _5 - _3;
    assign _7 = funct7;
    assign _22 = _7[0:0];
    assign _25 = _22 ? _24 : _23;
    assign _9 = funct3;
    always @* begin
        case (_9)
        0: _486 <= _25;
        1: _486 <= _123;
        2: _486 <= _134;
        3: _486 <= _137;
        4: _486 <= _138;
        5: _486 <= _483;
        6: _486 <= _484;
        default: _486 <= _485;
        endcase
    end

    /* aliases */

    /* output assignments */
    assign new_rd = _486;
    assign error = _21;

endmodule
